module andgate (a,b,c);
input a,b;
output c;
assign c=a&b;
endmodule 

module andgate_tb;


//test bench

module andgate_tb();
reg a,b;
wire c;
andgate OUT (.a(a),.b(b),.c(c));
initial begin
$monitor("a=%b b=%b c=%b",a,b,c);
a=0;
b=0;
#10
a=0;
b=1;
#10
a=1;
b=0;
#10
a=1;
b=1;
#10;
end 
endmodule 


